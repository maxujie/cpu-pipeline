module ALU(
  input [31:0] A,
  input [31:0] B,
  input [5:0] ALUFun,
  input Sign,
  output [31:0] Z
  );

endmodule
