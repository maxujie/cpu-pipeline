module CPU_Pipeline (
  input clk,
  input reset_b);

wire [63:0] IF_ID;














end module
